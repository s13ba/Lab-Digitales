`timescale 1ns / 1ps

module sumador(
    input  A,B

    );
endmodule
