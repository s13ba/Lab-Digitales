`timescale 1ns / 1ps
//Contador de N bits (por defecto 4)
//Pregunta 3.7 gu�a 2

module nbit_counter #(parameter N=4)(
     input  logic          clk, reset, PB_in,
     output logic [N-1:0]  count

    );
    
    always_ff @(posedge clk) begin //flip flop
    //se activa al pasar por el canto de subida del reloj
        if (reset) //si se�al reset es 1...
            count <= 'd0; //contador se reinicia
        else
            if (PB_in)
                count <= count+1; //sino, va sumando en cada canto positivo
            else
                count <= count;
    end
endmodule
